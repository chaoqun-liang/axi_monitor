// Copyright 2023 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Authors:
// - Chaoqun Liang <chaoqun.liang@unibo.it>


// hmmmm, the one of xbar was not the best choice
// go with a simple one first
// one master and one slave first
