// take out queue from write and read